-- Loren Lugosch
-- ECSE 682 Project
-- 
-- rsqrt.vhd

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE work.parameters.all;

ENTITY rsqrt IS
	PORT(
		--clock : IN STD_LOGIC;
		--reset : IN STD_LOGIC;
		sum_2 : IN SIGNED(Q21_43.data_width-1 DOWNTO 0);
		w_rnorm : OUT SIGNED(Q11_21.data_width-1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE arch OF rsqrt IS

	SIGNAL a : SIGNED(Q11_21.data_width-1 DOWNTO 0);
	SIGNAL b : SIGNED(Q21_43.data_width-1 DOWNTO 0);
	SIGNAL c : SIGNED(Q21_43.data_width-1 DOWNTO 0);
	SIGNAL d : SIGNED(Q21_43.data_width-1 DOWNTO 0);
	SIGNAL e : SIGNED(Q21_43.data_width-1 DOWNTO 0);
	SIGNAL f : SIGNED(Q21_43.data_width-1 DOWNTO 0);

BEGIN

	PROCESS(sum_2)
	BEGIN

		IF ((sum_2 >=    "0000000000000000000000000000000000000000000000000000000000000000") AND (sum_2 < "0000000000000000101000000000000000000000000000000000000000000000")) 	THEN a <= "11111111111111110010000100111010"; b <= "0000000000000000000001010101001010001000110011100111000000111010"; e <= sum_2;
		ELSIF ((sum_2 >= "0000000000000000101000000000000000000000000000000000000000000000") AND (sum_2 < "0000000000000001010000000000000000000000000000000000000000000000")) 	THEN a <= "11111111111111111110010111011010"; b <= "0000000000000000000000100100000000011010001101101110001011101011"; e <= sum_2;
		ELSIF ((sum_2 >= "0000000000000001010000000000000000000000000000000000000000000000") AND (sum_2 < "0000000000000010010110000000000000000000000000000000000000000000")) 	THEN a <= "11111111111111111111011000111110"; b <= "0000000000000000000000011001110111100110100110101101010000101100"; e <= sum_2;
		ELSIF ((sum_2 >= "0000000000000010010110000000000000000000000000000000000000000000") AND (sum_2 < "0000000000000100101100000000000000000000000000000000000000000000")) 	THEN a <= "11111111111111111111110001101010"; b <= "0000000000000000000000010010100011110101110000101000111101011100"; e <= sum_2;
		ELSIF ((sum_2 >= "0000000000000100101100000000000000000000000000000000000000000000") AND (sum_2 < "0000000000000111110100000000000000000000000000000000000000000000")) 	THEN a <= "11111111111111111111111010000101"; b <= "0000000000000000000000001101110000101000111101011100001010001111"; e <= sum_2;
		ELSIF ((sum_2 >= "0000000000000111110100000000000000000000000000000000000000000000") AND (sum_2 < "0000000000001111101000000000000000000000000000000000000000000000")) 	THEN a <= "11111111111111111111111101101010"; b <= "0000000000000000000000001010001010011100011101111001101001101011"; e <= sum_2;
		ELSIF ((sum_2 >= "0000000000001111101000000000000000000000000000000000000000000000") AND (sum_2 < "0000000000011111010000000000000000000000000000000000000000000000")) 	THEN a <= "11111111111111111111111001010110"; b <= "0000000000000000000000000111001011100100100011101000101001110001"; e <= sum_2 srl 3;
		ELSE																																										 a <= "11111111111111111111111101101010"; b <= "0000000000000000000000000101000101001110001110111100110100110101"; e <= sum_2 srl 3;
		END IF;

	END PROCESS;

	--return (Q11_21)((multiply_Q11_21_by_Q11_21((Q11_21)(input >> 22),a) + b) >> 22);

	f <= (e srl 22);
	c <= ((a * f(Q11_21.data_width-1 DOWNTO 0)) sll 1) + b;
	d <= c srl 22;
	w_rnorm <= d(Q11_21.data_width-1 DOWNTO 0);

END arch;