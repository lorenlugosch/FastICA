-- Loren Lugosch
-- ECSE 682 Project
-- 
-- sech2.vhd

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE work.parameters.all;

ENTITY sech2 IS
	PORT(
		--clock : IN STD_LOGIC;
		--reset : IN STD_LOGIC;
		p1 : IN SIGNED(Q11_21.data_width-1 DOWNTO 0);
		sp : OUT SIGNED(Q11_21.data_width-1 DOWNTO 0)
	);
END ENTITY;

ARCHITECTURE arch OF sech2 IS
 
	SIGNAL a : SIGNED(Q11_21.data_width-1 DOWNTO 0);
	SIGNAL b : SIGNED(Q21_43.data_width-1 DOWNTO 0);
	SIGNAL c : SIGNED(Q21_43.data_width-1 DOWNTO 0);
	SIGNAL d : SIGNED(Q21_43.data_width-1 DOWNTO 0);

BEGIN

	PROCESS(p1)
	BEGIN

		IF    (p1 < "11111111101000000000000000000000") 													THEN a <= "00000000000000000001111110110011"; b <= "0000000000000000000000000010010010101000110000010101010011001001";
		ELSIF ((p1 >= "11111111101000000000000000000000") AND (p1 < "11111111110000000000000000000000")) 	THEN a <= "00000000000000011100111000101001"; b <= "0000000000000000000000010110000001110101111101101111110100100001";
		ELSIF ((p1 >= "11111111110000000000000000000000") AND (p1 < "11111111110100000000000000000000")) 	THEN a <= "00000000000001101101101001010001"; b <= "0000000000000000000000111111000011011000010001001101000000010011";
		ELSIF ((p1 >= "11111111110100000000000000000000") AND (p1 < "11111111111000000000000000000000")) 	THEN a <= "00000000000011110001010000100010"; b <= "0000000000000000000001110000001010101001100100110000101111100000";
		ELSIF ((p1 >= "11111111111000000000000000000000") AND (p1 < "11111111111100000000000000000000")) 	THEN a <= "00000000000101111010111101101010"; b <= "0000000000000000000010010011101111001101001101011010100001011000";
		ELSIF ((p1 >= "11111111111100000000000000000000") AND (p1 < "11111111111110011001100110011001")) 	THEN a <= "00000000000100110010100001011001"; b <= "0000000000000000000010001011110000000001101000110110111000101110";
		ELSIF ((p1 >= "11111111111110011001100110011001") AND (p1 < "00000000000000000000000000000000")) 	THEN a <= "00000000000001101101111001000111"; b <= "0000000000000000000010000001000010010110101110111001100011000111";	
		ELSIF ((p1 >= "00000000000000000000000000000000") AND (p1 < "00000000000001100110011001100110")) 	THEN a <= "11111111111110010010000110111001"; b <= "0000000000000000000010000001000010010110101110111001100011000111";
		ELSIF ((p1 >= "00000000000001100110011001100110") AND (p1 < "00000000000100000000000000000000")) 	THEN a <= "11111111111011001101011110100111"; b <= "0000000000000000000010001011110000000001101000110110111000101110";
		ELSIF ((p1 >= "00000000000100000000000000000000") AND (p1 < "00000000001000000000000000000000"))	THEN a <= "11111111111010000101000010010110"; b <= "0000000000000000000010010011101111001101001101011010100001011000";
		ELSIF ((p1 >= "00000000001000000000000000000000") AND (p1 < "00000000001100000000000000000000")) 	THEN a <= "11111111111100001110101111011110"; b <= "0000000000000000000001110000001010101001100100110000101111100000";
		ELSIF ((p1 >= "00000000001100000000000000000000") AND (p1 < "00000000010000000000000000000000")) 	THEN a <= "11111111111110010010010110101111"; b <= "0000000000000000000000111111000011011000010001001101000000010011";
		ELSIF ((p1 >= "00000000010000000000000000000000") AND (p1 < "00000000011000000000000000000000")) 	THEN a <= "11111111111111100011000111010111"; b <= "0000000000000000000000010110000001110101111101101111110100100001";
		ELSE																									 a <= "11111111111111111110000001001101"; b <= "0000000000000000000000000010010010101000110000010101010011001001";
		END IF;

	END PROCESS;

	c <= ((a * p1) sll 1) + b;
	d <= c srl 22;
	sp <= d(Q11_21.data_width-1 DOWNTO 0);

END arch;